`ifndef sys_array_defines
    `define sys_array_defines
        enum {simple, load} sys_array_cell_types;
`endif
